`define I_CACHE_INDEX   12
`define D_CACHE_INDEX   11

`define PLL_FREQ        clk_pll
`define I_CACHE_INDEX   6
`define D_CACHE_INDEX   6

`define PLL_FREQ        clk_pll
`define I_CACHE_INDEX   8
`define D_CACHE_INDEX   8

`define PLL_FREQ        clk_pll_80
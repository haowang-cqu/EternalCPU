`define I_CACHE_INDEX   5
`define D_CACHE_INDEX   5
`define I_CACHE_WRD_INDEX 4 
`define D_CACHE_WRD_INDEX 4

`define PLL_FREQ        clk_pll
// Cache Config
`define I_CACHE_INDEX   4
`define D_CACHE_INDEX   4
`define I_CACHE_WRD_INDEX 4 
`define D_CACHE_WRD_INDEX 4
// PLL Config
`define PLL_FREQ        clk_pll_85
// TLB Config
`define ENABLE_TLB      1
`define TLB_WIDTH       5
`define TLB_LINE        (1<<`TLB_WIDTH)
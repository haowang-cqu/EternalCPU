// Cache Config
`define I_CACHE_INDEX   12
`define D_CACHE_INDEX   11
// PLL Config
`define PLL_FREQ        clk_pll
// TLB Config
`define ENABLE_TLB      0
`define TLB_WIDTH       5
`define TLB_LINE        (1<<`TLB_WIDTH)
`timescale 1ns / 1ps

`include "defines.vh"
module branch_controller(
	input  wire [31:0] rdata1_i,
	input  wire [31:0] rdata2_i,
	input  wire [5:0]  id_op_i,
	input  wire [4:0]  id_rt_i,
	output reg         id_equal_o
    );
	always@(*) begin
		case(id_op_i)
			`BEQ,  `BEQL : id_equal_o <= (rdata1_i == rdata2_i) ? 1 : 0;
			`BNE,  `BNEL : id_equal_o <= (rdata1_i == rdata2_i) ? 0 : 1;
			`BGTZ, `BGTZL: id_equal_o <= (rdata1_i[31] == 0 && rdata1_i != 32'b0) ? 1: 0;
			`BLEZ, `BLEZL: id_equal_o <= (rdata1_i[31] == 1 || rdata1_i == 32'b0) ? 1: 0;
			`REGIMM_INST:case(id_rt_i)
							`BLTZ,   `BLTZL  : id_equal_o <= (rdata1_i[31] == 1) ? 1: 0;
							`BLTZAL, `BLTZALL: id_equal_o <= (rdata1_i[31] == 1) ? 1: 0;
							`BGEZ,   `BGEZL  : id_equal_o <= (rdata1_i[31] == 0) ? 1: 0;
							`BGEZAL, `BGEZALL: id_equal_o <= (rdata1_i[31] == 0) ? 1: 0;
							default:id_equal_o <= 0;
						 endcase
			default:id_equal_o<=0;
		endcase
	end
endmodule
